`ifndef DEFINES_H
  `define DEFINES_H

  `define NUMNODES 4
  `define PORT_RING 18244
  `define PORT_CROSSBAR 18241
  `define PORT_MESH 18242
  `define PORT_BUS 18243
  `define CLOCK_RATIO 8
`endif