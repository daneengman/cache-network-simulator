`define VERBOSE