`default_nettype none

module ring (
  input clk, rst_l
);

endmodule: ring