`default_nettype none

module bus (
  input clk, rst_l
);

endmodule: bus