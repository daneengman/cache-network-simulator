`default_nettype none

module top();

  logic clk, rst_l;

  ring dut(.*);

  

endmodule: top